// Register file

module register_file(output reg [31:0] out, input [31:0] in, input enable, Clr, Clk); // still missing some arguments