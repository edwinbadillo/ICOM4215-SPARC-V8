// 32 bit 2x1 Multiplexer
module mux_2x1 (output reg [31: 0]Y, input S, [31: 0]I0, [31: 0]I1); 
always @ (S, I0, I1) 
if (S) Y = I1; 
else Y = I0; 
endmodule

// 32 bit 4x1 Multiplexer
module mux_4x1 (output reg [31: 0]Y, input [1:0]S, [31: 0]I0, [31:0]I1, [31:0]I2, [31:0]I3); 
always @ (S, I0, I1, I2, I3) 
case(S)
2'b00: Y = I0; 
2'b01: Y = I1; 
2'b10: Y = I2; 
2'b11: Y = I3; 
endcase
endmodule


// 32 bit 8x1 Multiplexer
module mux_8x1 (output reg [31: 0]Y, input [3:0]S, [31: 0]I0, [31:0]I1, [31:0]I2, [31:0]I3, [31:0]I4, [31:0]I5, [31:0]I6, [31:0]I7, [31:0]I8); 
always @ (S, I0, I1, I2, I3, I4, I5, I6, I7) 
case(S)
3'b000: Y = I0; 
3'b001: Y = I1; 
3'b010: Y = I2; 
3'b011: Y = I3; 
3'b100: Y = I4; 
3'b101: Y = I5; 
3'b110: Y = I6; 
3'b111: Y = I7;

endcase
endmodule

// 32 bit 64x1 Multiplexer
module mux_64x1 (output reg [31: 0]Y, input [5:0]S, reg[31:0] I[0:63]); 
always @ (S, I) 
case(S)
6'b000000: Y = I[000000];
6'b000001: Y = I[000001];
6'b000010: Y = I[000010];
6'b000011: Y = I[000011];
6'b000100: Y = I[000100];
6'b000101: Y = I[000101];
6'b000110: Y = I[000110];
6'b000111: Y = I[000111];
6'b001000: Y = I[001000];
6'b001001: Y = I[001001];
6'b001010: Y = I[001010];
6'b001011: Y = I[001011];
6'b001100: Y = I[001100];
6'b001101: Y = I[001101];
6'b001110: Y = I[001110];
6'b001111: Y = I[001111];
6'b010000: Y = I[010000];
6'b010001: Y = I[010001];
6'b010010: Y = I[010010];
6'b010011: Y = I[010011];
6'b010100: Y = I[010100];
6'b010101: Y = I[010101];
6'b010110: Y = I[010110];
6'b010111: Y = I[010111];
6'b011000: Y = I[011000];
6'b011001: Y = I[011001];
6'b011010: Y = I[011010];
6'b011011: Y = I[011011];
6'b011100: Y = I[011100];
6'b011101: Y = I[011101];
6'b011110: Y = I[011110];
6'b011111: Y = I[011111];
6'b100000: Y = I[100000];
6'b100001: Y = I[100001];
6'b100010: Y = I[100010];
6'b100011: Y = I[100011];
6'b100100: Y = I[100100];
6'b100101: Y = I[100101];
6'b100110: Y = I[100110];
6'b100111: Y = I[100111];
6'b101000: Y = I[101000];
6'b101001: Y = I[101001];
6'b101010: Y = I[101010];
6'b101011: Y = I[101011];
6'b101100: Y = I[101100];
6'b101101: Y = I[101101];
6'b101110: Y = I[101110];
6'b101111: Y = I[101111];
6'b110000: Y = I[110000];
6'b110001: Y = I[110001];
6'b110010: Y = I[110010];
6'b110011: Y = I[110011];
6'b110100: Y = I[110100];
6'b110101: Y = I[110101];
6'b110110: Y = I[110110];
6'b110111: Y = I[110111];
6'b111000: Y = I[111000];
6'b111001: Y = I[111001];
6'b111010: Y = I[111010];
6'b111011: Y = I[111011];
6'b111100: Y = I[111100];
6'b111101: Y = I[111101];
6'b111110: Y = I[111110];
6'b111111: Y = I[111111];
endcase
endmodule
