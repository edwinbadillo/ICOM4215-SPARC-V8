// Register file

module register_file(output reg [31:0] out, input [31:0] in, input enable, Clr, Clk, current_window); // still missing some arguments


decoder_2x4()



//DFF d[15:0] (clk, DFF_i, DFF_o);


endmodule
